//-----------------------------------------------------------------------------
// Copyright 2021 Andrea Miele
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//-----------------------------------------------------------------------------

// qSelPLAPos.sv
// Non-negative only PLA for Radix-4 SRT quotient selection 
// -2/3y <= r <= 2/3 y
// follows table in H&P 5th edition, appendix J, page 57

module qSelPLAPos
(
    input logic [4 : 0] r5,
    input logic [3 : 0] y4,
    output logic [1 : 0] q2 // magnitude of quotient digit 
);

always_comb
begin

    case ({y4, r5})
        // 8 0: 0
        {4'h8, 5'h0}: q2 = 2'b00;
        // 8 1: 0
        {4'h8, 5'h1}: q2 = 2'b00;
        // 8 2: 1
        {4'h8, 5'h2}: q2 = 2'b01;
        // 8 3: 1
        {4'h8, 5'h3}: q2 = 2'b01;
        // 8 4: 1
        {4'h8, 5'h4}: q2 = 2'b01;
        // 8 5: 1
        {4'h8, 5'h5}: q2 = 2'b01;
        // 8 6: 2
        {4'h8, 5'h6}: q2 = 2'b10;
        // 8 7: 2
        {4'h8, 5'h7}: q2 = 2'b10;
        // 8 8: 2
        {4'h8, 5'h8}: q2 = 2'b10;
        // 8 9: 2
        {4'h8, 5'h9}: q2 = 2'b10;
        // 8 10: 2
        {4'h8, 5'ha}: q2 = 2'b10;
        // 8 11: 2
        {4'h8, 5'hb}: q2 = 2'b10;
        // 9 0: 0
        {4'h9, 5'h0}: q2 = 2'b00;
        // 9 1: 0
        {4'h9, 5'h1}: q2 = 2'b00;
        // 9 2: 0
        {4'h9, 5'h2}: q2 = 2'b00;
        // 9 3: 1
        {4'h9, 5'h3}: q2 = 2'b01;
        // 9 4: 1
        {4'h9, 5'h4}: q2 = 2'b01;
        // 9 5: 1
        {4'h9, 5'h5}: q2 = 2'b01;
        // 9 6: 1
        {4'h9, 5'h6}: q2 = 2'b01;
        // 9 7: 2
        {4'h9, 5'h7}: q2 = 2'b10;
        // 9 8: 2
        {4'h9, 5'h8}: q2 = 2'b10;
        // 9 9: 2
        {4'h9, 5'h9}: q2 = 2'b10;
        // 9 10: 2
        {4'h9, 5'ha}: q2 = 2'b10;
        // 9 11: 2
        {4'h9, 5'hb}: q2 = 2'b10;
        // 9 12: 2
        {4'h9, 5'hc}: q2 = 2'b10;
        // 9 13: 2
        {4'h9, 5'hd}: q2 = 2'b10;
        // 10 0: 0
        {4'ha, 5'h0}: q2 = 2'b00;
        // 10 1: 0
        {4'ha, 5'h1}: q2 = 2'b00;
        // 10 2: 0
        {4'ha, 5'h2}: q2 = 2'b00;
        // 10 3: 1
        {4'ha, 5'h3}: q2 = 2'b01;
        // 10 4: 1
        {4'ha, 5'h4}: q2 = 2'b01;
        // 10 5: 1
        {4'ha, 5'h5}: q2 = 2'b01;
        // 10 6: 1
        {4'ha, 5'h6}: q2 = 2'b01;
        // 10 7: 1
        {4'ha, 5'h7}: q2 = 2'b01;
        // 10 8: 2
        {4'ha, 5'h8}: q2 = 2'b10;
        // 10 9: 2
        {4'ha, 5'h9}: q2 = 2'b10;
        // 10 10: 2
        {4'ha, 5'ha}: q2 = 2'b10;
        // 10 11: 2
        {4'ha, 5'hb}: q2 = 2'b10;
        // 10 12: 2
        {4'ha, 5'hc}: q2 = 2'b10;
        // 10 13: 2
        {4'ha, 5'hd}: q2 = 2'b10;
        // 10 14: 2
        {4'ha, 5'he}: q2 = 2'b10;
        // 11 0: 0
        {4'hb, 5'h0}: q2 = 2'b00;
        // 11 1: 0
        {4'hb, 5'h1}: q2 = 2'b00;
        // 11 2: 0
        {4'hb, 5'h2}: q2 = 2'b00;
        // 11 3: 1
        {4'hb, 5'h3}: q2 = 2'b01;
        // 11 4: 1
        {4'hb, 5'h4}: q2 = 2'b01;
        // 11 5: 1
        {4'hb, 5'h5}: q2 = 2'b01;
        // 11 6: 1
        {4'hb, 5'h6}: q2 = 2'b01;
        // 11 7: 1
        {4'hb, 5'h7}: q2 = 2'b01;
        // 11 8: 1
        {4'hb, 5'h8}: q2 = 2'b01;
        // 11 9: 2
        {4'hb, 5'h9}: q2 = 2'b10;
        // 11 10: 2
        {4'hb, 5'ha}: q2 = 2'b10;
        // 11 11: 2
        {4'hb, 5'hb}: q2 = 2'b10;
        // 11 12: 2
        {4'hb, 5'hc}: q2 = 2'b10;
        // 11 13: 2
        {4'hb, 5'hd}: q2 = 2'b10;
        // 11 14: 2
        {4'hb, 5'he}: q2 = 2'b10;
        // 11 15: 2
        {4'hb, 5'hf}: q2 = 2'b10;
        // 12 0: 0
        {4'hc, 5'h0}: q2 = 2'b00;
        // 12 1: 0
        {4'hc, 5'h1}: q2 = 2'b00;
        // 12 2: 0
        {4'hc, 5'h2}: q2 = 2'b00;
        // 12 3: 0
        {4'hc, 5'h3}: q2 = 2'b00;
        // 12 4: 1
        {4'hc, 5'h4}: q2 = 2'b01;
        // 12 5: 1
        {4'hc, 5'h5}: q2 = 2'b01;
        // 12 6: 1
        {4'hc, 5'h6}: q2 = 2'b01;
        // 12 7: 1
        {4'hc, 5'h7}: q2 = 2'b01;
        // 12 8: 1
        {4'hc, 5'h8}: q2 = 2'b01;
        // 12 9: 1
        {4'hc, 5'h9}: q2 = 2'b01;
        // 12 10: 2
        {4'hc, 5'ha}: q2 = 2'b10;
        // 12 11: 2
        {4'hc, 5'hb}: q2 = 2'b10;
        // 12 12: 2
        {4'hc, 5'hc}: q2 = 2'b10;
        // 12 13: 2
        {4'hc, 5'hd}: q2 = 2'b10;
        // 12 14: 2
        {4'hc, 5'he}: q2 = 2'b10;
        // 12 15: 2
        {4'hc, 5'hf}: q2 = 2'b10;
        // 12 16: 2
        {4'hc, 5'h10}: q2 = 2'b10;
        // 12 17: 2
        {4'hc, 5'h11}: q2 = 2'b10;
        // 13 0: 0
        {4'hd, 5'h0}: q2 = 2'b00;
        // 13 1: 0
        {4'hd, 5'h1}: q2 = 2'b00;
        // 13 2: 0
        {4'hd, 5'h2}: q2 = 2'b00;
        // 13 3: 0
        {4'hd, 5'h3}: q2 = 2'b00;
        // 13 4: 1
        {4'hd, 5'h4}: q2 = 2'b01;
        // 13 5: 1
        {4'hd, 5'h5}: q2 = 2'b01;
        // 13 6: 1
        {4'hd, 5'h6}: q2 = 2'b01;
        // 13 7: 1
        {4'hd, 5'h7}: q2 = 2'b01;
        // 13 8: 1
        {4'hd, 5'h8}: q2 = 2'b01;
        // 13 9: 1
        {4'hd, 5'h9}: q2 = 2'b01;
        // 13 10: 2
        {4'hd, 5'ha}: q2 = 2'b10;
        // 13 11: 2
        {4'hd, 5'hb}: q2 = 2'b10;
        // 13 12: 2
        {4'hd, 5'hc}: q2 = 2'b10;
        // 13 13: 2
        {4'hd, 5'hd}: q2 = 2'b10;
        // 13 14: 2
        {4'hd, 5'he}: q2 = 2'b10;
        // 13 15: 2
        {4'hd, 5'hf}: q2 = 2'b10;
        // 13 16: 2
        {4'hd, 5'h10}: q2 = 2'b10;
        // 13 17: 2
        {4'hd, 5'h11}: q2 = 2'b10;
        // 13 18: 2
        {4'hd, 5'h12}: q2 = 2'b10;
        // 14 0: 0
        {4'he, 5'h0}: q2 = 2'b00;
        // 14 1: 0
        {4'he, 5'h1}: q2 = 2'b00;
        // 14 2: 0
        {4'he, 5'h2}: q2 = 2'b00;
        // 14 3: 0
        {4'he, 5'h3}: q2 = 2'b00;
        // 14 4: 1
        {4'he, 5'h4}: q2 = 2'b01;
        // 14 5: 1
        {4'he, 5'h5}: q2 = 2'b01;
        // 14 6: 1
        {4'he, 5'h6}: q2 = 2'b01;
        // 14 7: 1
        {4'he, 5'h7}: q2 = 2'b01;
        // 14 8: 1
        {4'he, 5'h8}: q2 = 2'b01;
        // 14 9: 1
        {4'he, 5'h9}: q2 = 2'b01;
        // 14 10: 1
        {4'he, 5'ha}: q2 = 2'b01;
        // 14 11: 2
        {4'he, 5'hb}: q2 = 2'b10;
        // 14 12: 2
        {4'he, 5'hc}: q2 = 2'b10;
        // 14 13: 2
        {4'he, 5'hd}: q2 = 2'b10;
        // 14 14: 2
        {4'he, 5'he}: q2 = 2'b10;
        // 14 15: 2
        {4'he, 5'hf}: q2 = 2'b10;
        // 14 16: 2
        {4'he, 5'h10}: q2 = 2'b10;
        // 14 17: 2
        {4'he, 5'h11}: q2 = 2'b10;
        // 14 18: 2
        {4'he, 5'h12}: q2 = 2'b10;
        // 14 19: 2
        {4'he, 5'h13}: q2 = 2'b10;
        // 15 0: 0
        {4'hf, 5'h0}: q2 = 2'b00;
        // 15 1: 0
        {4'hf, 5'h1}: q2 = 2'b00;
        // 15 2: 0
        {4'hf, 5'h2}: q2 = 2'b00;
        // 15 3: 0
        {4'hf, 5'h3}: q2 = 2'b00;
        // 15 4: 0
        {4'hf, 5'h4}: q2 = 2'b00;
        // 15 5: 1
        {4'hf, 5'h5}: q2 = 2'b01;
        // 15 6: 1
        {4'hf, 5'h6}: q2 = 2'b01;
        // 15 7: 1
        {4'hf, 5'h7}: q2 = 2'b01;
        // 15 8: 1
        {4'hf, 5'h8}: q2 = 2'b01;
        // 15 9: 1
        {4'hf, 5'h9}: q2 = 2'b01;
        // 15 10: 1
        {4'hf, 5'ha}: q2 = 2'b01;
        // 15 11: 1
        {4'hf, 5'hb}: q2 = 2'b01;
        // 15 12: 2
        {4'hf, 5'hc}: q2 = 2'b10;
        // 15 13: 2
        {4'hf, 5'hd}: q2 = 2'b10;
        // 15 14: 2
        {4'hf, 5'he}: q2 = 2'b10;
        // 15 15: 2
        {4'hf, 5'hf}: q2 = 2'b10;
        // 15 16: 2
        {4'hf, 5'h10}: q2 = 2'b10;
        // 15 17: 2
        {4'hf, 5'h11}: q2 = 2'b10;
        // 15 18: 2
        {4'hf, 5'h12}: q2 = 2'b10;
        // 15 19: 2
        {4'hf, 5'h13}: q2 = 2'b10;
        // 15 20: 2
        {4'hf, 5'h14}: q2 = 2'b10;
        // 15 21: 2
        {4'hf, 5'h15}: q2 = 2'b10;
		  
		  default:       q2 = 2'b00;

    endcase
end
endmodule
